//===========================================================================
// Module name: key_test.v
// ����: ��⿪�����ϵ��ĸ�����KEY1~KEY4, ����⵽��������ʱ,��Ӧ��LED�Ʒ�ת
//===========================================================================
`timescale 1ns / 1ps
module key_test  (
							clk,              // ������������ʱ��: 50Mhz
							rst_n,            // �����������븴λ����
							key_in,           // ���밴���ź�(KEY1~KEY4)
							out           // ���LED��,���ڿ��ƿ��������ĸ�LED(LED1~LED4)
						);

//===========================================================================
// PORT declarations
//===========================================================================						
input        clk; 
input        rst_n;
input  [5:0] key_in;
output [5:0] out;

//�Ĵ�������
reg [19:0] count;
reg [5:0] key_scan; //����ɨ��ֵKEY

//===========================================================================
// ��������ֵ��20msɨ��һ��,����Ƶ��С�ڰ���ë��Ƶ�ʣ��൱���˳����˸�Ƶë���źš�
//===========================================================================
always @(posedge clk or negedge rst_n)     //���ʱ�ӵ������غ͸�λ���½���
begin
   if(!rst_n)                //��λ�źŵ���Ч
      count <= 20'd0;        //��������0
   else
      begin
         if(count ==20'd999_999)   //20msɨ��һ�ΰ���,20ms����(50M/50-1=999_999)
            begin
               count <= 20'b0;     //�������Ƶ�20ms������������
               key_scan <= key_in; //�������������ƽ
            end
         else
            count <= count + 20'b1; //��������1
     end
end
//===========================================================================
// �����ź�����һ��ʱ�ӽ���
//===========================================================================
reg [5:0] key_scan_r;
always @(posedge clk)
    key_scan_r <= key_scan;       
    
wire [5:0] flag_key = key_scan_r[5:0] & (~key_scan[5:0]);  //����⵽�������½��ر仯ʱ������ð��������£�������Ч 
assign out = flag_key;
//===========================================================================

endmodule

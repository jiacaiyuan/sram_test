module  SRAM_SOC
	(
		////////////////////	Clock Input	 	////////////////////	 
		
		CLOCK_50,						//	On Board 50 MHz
		////////////////////	Push Button		////////////////////
		KEY,							//	Pushbutton[3:0]
		////////////////////////	LED		////////////////////////
		LEDG,							//	LED Green[8:0]
		////////////////////////	IP_INTERFACE	///////////////
		s_clk,
		s_cen,
		s_oen,
		s_wen,
		s_addr,
		s_ddata,
		s_qdata,
		/////////////////////	SDRAM Interface		////////////////
		DRAM_DQ,						//	SDRAM Data bus 16 Bits
		DRAM_ADDR,						//	SDRAM Address bus 12 Bits
		DRAM_LDQM,						//	SDRAM Low-byte Data Mask 
		DRAM_UDQM,						//	SDRAM High-byte Data Mask
		DRAM_WE_N,						//	SDRAM Write Enable
		DRAM_CAS_N,						//	SDRAM Column Address Strobe
		DRAM_RAS_N,						//	SDRAM Row Address Strobe
		DRAM_CS_N,						//	SDRAM Chip Select
		DRAM_BA_0,						//	SDRAM Bank Address 0
		DRAM_BA_1,						//	SDRAM Bank Address 1
		DRAM_CLK,						//	SDRAM Clock
		DRAM_CKE,						//	SDRAM Clock Enable
		////////////	Ethernet Interface	////////////////////////
		ENET_DATA,						//	DM9000A DATA bus 16Bits
		ENET_CMD,						//	DM9000A Command/Data Select, 0 = Command, 1 = Data
		ENET_CS_N,						//	DM9000A Chip Select
		ENET_WR_N,						//	DM9000A Write
		ENET_RD_N,						//	DM9000A Read
		ENET_RST_N,						//	DM9000A Reset
		ENET_INT,						//	DM9000A Interrupt
		ENET_CLK						//	DM9000A Clock 25 MHz
	
		
		////////////////////	GPIO	////////////////////////////
/*		GPIO_0,							//	GPIO Connection 0
		GPIO_1							//	GPIO Connection 1
*/
		
	);
	
	////////////////////////	Clock Input	 	////////////////////////

input			CLOCK_50;				//	On Board 50 MHz

////////////////////////	Push Button		////////////////////////
input	[3:0]	KEY;					//	Pushbutton[3:0]
////////////////////////	IP_INTERFACE		////////////////////////
output	s_clk;
output	s_cen;
output	s_oen;
output	s_wen;

input	[7:0]	s_qdata;	
output	[7:0]	s_ddata;
output	[9:0]	s_addr;
////////////////////////////	LED		////////////////////////////

output	[8:0]	LEDG;					//	LED Green[8:0]



///////////////////////		SDRAM Interface	////////////////////////
inout	[15:0]	DRAM_DQ;				//	SDRAM Data bus 16 Bits
output	[11:0]	DRAM_ADDR;				//	SDRAM Address bus 12 Bits
output			DRAM_LDQM;				//	SDRAM Low-byte Data Mask 
output			DRAM_UDQM;				//	SDRAM High-byte Data Mask
output			DRAM_WE_N;				//	SDRAM Write Enable
output			DRAM_CAS_N;				//	SDRAM Column Address Strobe
output			DRAM_RAS_N;				//	SDRAM Row Address Strobe
output			DRAM_CS_N;				//	SDRAM Chip Select
output			DRAM_BA_0;				//	SDRAM Bank Address 0
output			DRAM_BA_1;				//	SDRAM Bank Address 0
output			DRAM_CLK;				//	SDRAM Clock
output			DRAM_CKE;				//	SDRAM Clock Enable

////////////////	Ethernet Interface	////////////////////////////

inout	[15:0]	ENET_DATA;				//	DM9000A DATA bus 16Bits
output			ENET_CMD;				//	DM9000A Command/Data Select, 0 = Command, 1 = Data
output			ENET_CS_N;				//	DM9000A Chip Select
output			ENET_WR_N;				//	DM9000A Write
output			ENET_RD_N;				//	DM9000A Read
output			ENET_RST_N;				//	DM9000A Reset
input			ENET_INT;				//	DM9000A Interrupt

output			ENET_CLK;				//	DM9000A Clock 25 MHz







////////////////////////	GPIO	////////////////////////////////
//inout	[35:0]	GPIO_0;					//	GPIO Connection 0
//inout	[35:0]	GPIO_1;					//	GPIO Connection 1

wire	CPU_CLK;
wire	CPU_RESET;
wire	ip_clk;



Reset_Delay	delay1	(.iRST(KEY[0]),.iCLK(CLOCK_50),.oRESET(CPU_RESET));
SDRAM_PLL 	PLL1	(.inclk0(CLOCK_50),.c0(DRAM_CLK),.c1(CPU_CLK),.c2(ip_clk));
											
system0 	u0	(
				// 1) global signals:
                  .clk_cpu(CPU_CLK),
                  .clk_sdram(CLOCK_50),
                  .reset_n(CPU_RESET),
				 // the_avalon_wrapper_0
				  .clk_to_the_avalon_wrapper_0(ip_clk),
                  .led_0_from_the_avalon_wrapper_0(LEDG[0]),
                  .led_1_from_the_avalon_wrapper_0(LEDG[1]),
                  .led_2_from_the_avalon_wrapper_0(LEDG[2]),
                  .led_3_from_the_avalon_wrapper_0(LEDG[3]),
                  .s_addr_from_the_avalon_wrapper_0(s_addr),
                  .s_cen_from_the_avalon_wrapper_0(s_cen),
                  .s_clk_from_the_avalon_wrapper_0(s_clk),
                  .s_ddata_from_the_avalon_wrapper_0(s_ddata),
                  .s_oen_from_the_avalon_wrapper_0(s_oen),
                  .s_qdata_to_the_avalon_wrapper_0(s_qdata),
                  .s_wen_from_the_avalon_wrapper_0(s_wen),
				 
                 // the_sdram_0
                 .zs_addr_from_the_sdram(DRAM_ADDR),
                 .zs_ba_from_the_sdram({DRAM_BA_1,DRAM_BA_0}),
                 .zs_cas_n_from_the_sdram(DRAM_CAS_N),
                 .zs_cke_from_the_sdram(DRAM_CKE),
                 .zs_cs_n_from_the_sdram(DRAM_CS_N),
                 .zs_dq_to_and_from_the_sdram(DRAM_DQ),
                 .zs_dqm_from_the_sdram({DRAM_UDQM,DRAM_LDQM}),
                 .zs_ras_n_from_the_sdram(DRAM_RAS_N),
                 .zs_we_n_from_the_sdram(DRAM_WE_N),
					  
					 
				// the_dm9000a_0
                  .ENET_CLK_from_the_dm9000a_0(ENET_CLK),
                  .ENET_CMD_from_the_dm9000a_0(ENET_CMD),
                  .ENET_CS_N_from_the_dm9000a_0(ENET_CS_N),
                  .ENET_DATA_to_and_from_the_dm9000a_0(ENET_DATA),
                  .ENET_INT_to_the_dm9000a_0(ENET_INT),
                  .ENET_RD_N_from_the_dm9000a_0(ENET_RD_N),
                  .ENET_RST_N_from_the_dm9000a_0(ENET_RST_N),
                  .ENET_WR_N_from_the_dm9000a_0(ENET_WR_N),
                  .iOSC_50_to_the_dm9000a_0(CLOCK_50)
						
						
					
                );	
endmodule
